module RegFile();



endmodule
